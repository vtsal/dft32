library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity realcoeff32 is
    generic(SIZE: integer;
	        WIDTH: integer:=18);
	port(
        index 		: in  std_logic_vector(2*SIZE-1 downto 0);
        coeff 		: out std_logic_vector(WIDTH-1 downto 0)
    );
end realcoeff32;

ARCHITECTURE dataflow OF realcoeff32 IS

SIGNAL indx: INTEGER RANGE 0 TO (2**SIZE)*(2**SIZE)-1;
TYPE vector_array IS ARRAY (0 to (2**SIZE)*(2**SIZE)-1) OF STD_LOGIC_VECTOR(20-1 DOWNTO 0);
CONSTANT memory : vector_array := 
	(
--32 point coefficients
--Row 0
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
--Row 1
x"00400",
x"003ec",
x"003b2",
x"00353",
x"002d4",
x"00238",
x"0030f",
x"0031f",
x"00000",
x"3fce1",
x"3fcf1",
x"3fdc8",
x"3fd2c",
x"3fcad",
x"3fc4e",
x"3fc14",
x"3fc00",
x"3fc14",
x"3fc4e",
x"3fcad",
x"3fd2c",
x"3fdc8",
x"3fcf1",
x"3fce1",
x"00000",
x"0031f",
x"0030f",
x"00238",
x"002d4",
x"00353",
x"003b2",
x"003ec",
--Row 2
x"00400",
x"003b2",
x"002d4",
x"0030f",
x"00000",
x"3fcf1",
x"3fd2c",
x"3fc4e",
x"3fc00",
x"3fc4e",
x"3fd2c",
x"3fcf1",
x"00000",
x"0030f",
x"002d4",
x"003b2",
x"00400",
x"003b2",
x"002d4",
x"0030f",
x"00000",
x"3fcf1",
x"3fd2c",
x"3fc4e",
x"3fc00",
x"3fc4e",
x"3fd2c",
x"3fcf1",
x"00000",
x"0030f",
x"002d4",
x"003b2",
--Row 3
x"00400",
x"00353",
x"0030f",
x"3fce1",
x"3fd2c",
x"3fc14",
x"3fc4e",
x"3fdc8",
x"00000",
x"00238",
x"003b2",
x"003ec",
x"002d4",
x"0031f",
x"3fcf1",
x"3fcad",
x"3fc00",
x"3fcad",
x"3fcf1",
x"0031f",
x"002d4",
x"003ec",
x"003b2",
x"00238",
x"00000",
x"3fdc8",
x"3fc4e",
x"3fc14",
x"3fd2c",
x"3fce1",
x"0030f",
x"00353",
--Row 4
x"00400",
x"002d4",
x"00000",
x"3fd2c",
x"3fc00",
x"3fd2c",
x"00000",
x"002d4",
x"00400",
x"002d4",
x"00000",
x"3fd2c",
x"3fc00",
x"3fd2c",
x"00000",
x"002d4",
x"00400",
x"002d4",
x"00000",
x"3fd2c",
x"3fc00",
x"3fd2c",
x"00000",
x"002d4",
x"00400",
x"002d4",
x"00000",
x"3fd2c",
x"3fc00",
x"3fd2c",
x"00000",
x"002d4",
--Row 5
x"00400",
x"00238",
x"3fcf1",
x"3fc14",
x"3fd2c",
x"0031f",
x"003b2",
x"00353",
x"00000",
x"3fcad",
x"3fc4e",
x"3fce1",
x"002d4",
x"003ec",
x"0030f",
x"3fdc8",
x"3fc00",
x"3fdc8",
x"0030f",
x"003ec",
x"002d4",
x"3fce1",
x"3fc4e",
x"3fcad",
x"00000",
x"00353",
x"003b2",
x"0031f",
x"3fd2c",
x"3fc14",
x"3fcf1",
x"00238",
--Row 6
x"00400",
x"0030f",
x"3fd2c",
x"3fc4e",
x"00000",
x"003b2",
x"002d4",
x"3fcf1",
x"3fc00",
x"3fcf1",
x"002d4",
x"003b2",
x"00000",
x"3fc4e",
x"3fd2c",
x"0030f",
x"00400",
x"0030f",
x"3fd2c",
x"3fc4e",
x"00000",
x"003b2",
x"002d4",
x"3fcf1",
x"3fc00",
x"3fcf1",
x"002d4",
x"003b2",
x"00000",
x"3fc4e",
x"3fd2c",
x"0030f",
--Row 7
x"00400",
x"0031f",
x"3fc4e",
x"3fdc8",
x"002d4",
x"00353",
x"3fcf1",
x"3fc14",
x"00000",
x"003ec",
x"0030f",
x"3fcad",
x"3fd2c",
x"00238",
x"003b2",
x"3fce1",
x"3fc00",
x"3fce1",
x"003b2",
x"00238",
x"3fd2c",
x"3fcad",
x"0030f",
x"003ec",
x"00000",
x"3fc14",
x"3fcf1",
x"00353",
x"002d4",
x"3fdc8",
x"3fc4e",
x"0031f",
--Row 8
x"00400",
x"00000",
x"3fc00",
x"00000",
x"00400",
x"00000",
x"3fc00",
x"00000",
x"00400",
x"00000",
x"3fc00",
x"00000",
x"00400",
x"00000",
x"3fc00",
x"00000",
x"00400",
x"00000",
x"3fc00",
x"00000",
x"00400",
x"00000",
x"3fc00",
x"00000",
x"00400",
x"00000",
x"3fc00",
x"00000",
x"00400",
x"00000",
x"3fc00",
x"00000",
--Row 9
x"00400",
x"3fce1",
x"3fc4e",
x"00238",
x"002d4",
x"3fcad",
x"3fcf1",
x"003ec",
x"00000",
x"3fc14",
x"0030f",
x"00353",
x"3fd2c",
x"3fdc8",
x"003b2",
x"0031f",
x"3fc00",
x"0031f",
x"003b2",
x"3fdc8",
x"3fd2c",
x"00353",
x"0030f",
x"3fc14",
x"00000",
x"003ec",
x"3fcf1",
x"3fcad",
x"002d4",
x"00238",
x"3fc4e",
x"3fce1",
--Row 10
x"00400",
x"3fcf1",
x"3fd2c",
x"003b2",
x"00000",
x"3fc4e",
x"002d4",
x"0030f",
x"3fc00",
x"0030f",
x"002d4",
x"3fc4e",
x"00000",
x"003b2",
x"3fd2c",
x"3fcf1",
x"00400",
x"3fcf1",
x"3fd2c",
x"003b2",
x"00000",
x"3fc4e",
x"002d4",
x"0030f",
x"3fc00",
x"0030f",
x"002d4",
x"3fc4e",
x"00000",
x"003b2",
x"3fd2c",
x"3fcf1",
--Row 11
x"00400",
x"3fdc8",
x"3fcf1",
x"003ec",
x"3fd2c",
x"3fce1",
x"003b2",
x"3fcad",
x"00000",
x"00353",
x"3fc4e",
x"0031f",
x"002d4",
x"3fc14",
x"0030f",
x"00238",
x"3fc00",
x"00238",
x"0030f",
x"3fc14",
x"002d4",
x"0031f",
x"3fc4e",
x"00353",
x"00000",
x"3fcad",
x"003b2",
x"3fce1",
x"3fd2c",
x"003ec",
x"3fcf1",
x"3fdc8",
--Row 12
x"00400",
x"3fd2c",
x"00000",
x"002d4",
x"3fc00",
x"002d4",
x"00000",
x"3fd2c",
x"00400",
x"3fd2c",
x"00000",
x"002d4",
x"3fc00",
x"002d4",
x"00000",
x"3fd2c",
x"00400",
x"3fd2c",
x"00000",
x"002d4",
x"3fc00",
x"002d4",
x"00000",
x"3fd2c",
x"00400",
x"3fd2c",
x"00000",
x"002d4",
x"3fc00",
x"002d4",
x"00000",
x"3fd2c",
--Row 13
x"00400",
x"3fcad",
x"0030f",
x"0031f",
x"3fd2c",
x"003ec",
x"3fc4e",
x"00238",
x"00000",
x"3fdc8",
x"003b2",
x"3fc14",
x"002d4",
x"3fce1",
x"3fcf1",
x"00353",
x"3fc00",
x"00353",
x"3fcf1",
x"3fce1",
x"002d4",
x"3fc14",
x"003b2",
x"3fdc8",
x"00000",
x"00238",
x"3fc4e",
x"003ec",
x"3fd2c",
x"0031f",
x"0030f",
x"3fcad",
--Row 14
x"00400",
x"3fc4e",
x"002d4",
x"3fcf1",
x"00000",
x"0030f",
x"3fd2c",
x"003b2",
x"3fc00",
x"003b2",
x"3fd2c",
x"0030f",
x"00000",
x"3fcf1",
x"002d4",
x"3fc4e",
x"00400",
x"3fc4e",
x"002d4",
x"3fcf1",
x"00000",
x"0030f",
x"3fd2c",
x"003b2",
x"3fc00",
x"003b2",
x"3fd2c",
x"0030f",
x"00000",
x"3fcf1",
x"002d4",
x"3fc4e",
--Row 15
x"00400",
x"3fc14",
x"003b2",
x"3fcad",
x"002d4",
x"3fdc8",
x"0030f",
x"3fce1",
x"00000",
x"0031f",
x"3fcf1",
x"00238",
x"3fd2c",
x"00353",
x"3fc4e",
x"003ec",
x"3fc00",
x"003ec",
x"3fc4e",
x"00353",
x"3fd2c",
x"00238",
x"3fcf1",
x"0031f",
x"00000",
x"3fce1",
x"0030f",
x"3fdc8",
x"002d4",
x"3fcad",
x"003b2",
x"3fc14",
--Row 16
x"00400",
x"3fc00",
x"00400",
x"3fc00",
x"00400",
x"3fc00",
x"00400",
x"3fc00",
x"00400",
x"3fc00",
x"00400",
x"3fc00",
x"00400",
x"3fc00",
x"00400",
x"3fc00",
x"00400",
x"3fc00",
x"00400",
x"3fc00",
x"00400",
x"3fc00",
x"00400",
x"3fc00",
x"00400",
x"3fc00",
x"00400",
x"3fc00",
x"00400",
x"3fc00",
x"00400",
x"3fc00",
--Row 17
x"00400",
x"3fc14",
x"003b2",
x"3fcad",
x"002d4",
x"3fdc8",
x"0030f",
x"3fce1",
x"00000",
x"0031f",
x"3fcf1",
x"00238",
x"3fd2c",
x"00353",
x"3fc4e",
x"003ec",
x"3fc00",
x"003ec",
x"3fc4e",
x"00353",
x"3fd2c",
x"00238",
x"3fcf1",
x"0031f",
x"00000",
x"3fce1",
x"0030f",
x"3fdc8",
x"002d4",
x"3fcad",
x"003b2",
x"3fc14",
--Row 18
x"00400",
x"3fc4e",
x"002d4",
x"3fcf1",
x"00000",
x"0030f",
x"3fd2c",
x"003b2",
x"3fc00",
x"003b2",
x"3fd2c",
x"0030f",
x"00000",
x"3fcf1",
x"002d4",
x"3fc4e",
x"00400",
x"3fc4e",
x"002d4",
x"3fcf1",
x"00000",
x"0030f",
x"3fd2c",
x"003b2",
x"3fc00",
x"003b2",
x"3fd2c",
x"0030f",
x"00000",
x"3fcf1",
x"002d4",
x"3fc4e",
--Row 19
x"00400",
x"3fcad",
x"0030f",
x"0031f",
x"3fd2c",
x"003ec",
x"3fc4e",
x"00238",
x"00000",
x"3fdc8",
x"003b2",
x"3fc14",
x"002d4",
x"3fce1",
x"3fcf1",
x"00353",
x"3fc00",
x"00353",
x"3fcf1",
x"3fce1",
x"002d4",
x"3fc14",
x"003b2",
x"3fdc8",
x"00000",
x"00238",
x"3fc4e",
x"003ec",
x"3fd2c",
x"0031f",
x"0030f",
x"3fcad",
--Row 20
x"00400",
x"3fd2c",
x"00000",
x"002d4",
x"3fc00",
x"002d4",
x"00000",
x"3fd2c",
x"00400",
x"3fd2c",
x"00000",
x"002d4",
x"3fc00",
x"002d4",
x"00000",
x"3fd2c",
x"00400",
x"3fd2c",
x"00000",
x"002d4",
x"3fc00",
x"002d4",
x"00000",
x"3fd2c",
x"00400",
x"3fd2c",
x"00000",
x"002d4",
x"3fc00",
x"002d4",
x"00000",
x"3fd2c",
--Row 21
x"00400",
x"3fdc8",
x"3fcf1",
x"003ec",
x"3fd2c",
x"3fce1",
x"003b2",
x"3fcad",
x"00000",
x"00353",
x"3fc4e",
x"0031f",
x"002d4",
x"3fc14",
x"0030f",
x"00238",
x"3fc00",
x"00238",
x"0030f",
x"3fc14",
x"002d4",
x"0031f",
x"3fc4e",
x"00353",
x"00000",
x"3fcad",
x"003b2",
x"3fce1",
x"3fd2c",
x"003ec",
x"3fcf1",
x"3fdc8",
--Row 22
x"00400",
x"3fcf1",
x"3fd2c",
x"003b2",
x"00000",
x"3fc4e",
x"002d4",
x"0030f",
x"3fc00",
x"0030f",
x"002d4",
x"3fc4e",
x"00000",
x"003b2",
x"3fd2c",
x"3fcf1",
x"00400",
x"3fcf1",
x"3fd2c",
x"003b2",
x"00000",
x"3fc4e",
x"002d4",
x"0030f",
x"3fc00",
x"0030f",
x"002d4",
x"3fc4e",
x"00000",
x"003b2",
x"3fd2c",
x"3fcf1",
--Row 23
x"00400",
x"3fce1",
x"3fc4e",
x"00238",
x"002d4",
x"3fcad",
x"3fcf1",
x"003ec",
x"00000",
x"3fc14",
x"0030f",
x"00353",
x"3fd2c",
x"3fdc8",
x"003b2",
x"0031f",
x"3fc00",
x"0031f",
x"003b2",
x"3fdc8",
x"3fd2c",
x"00353",
x"0030f",
x"3fc14",
x"00000",
x"003ec",
x"3fcf1",
x"3fcad",
x"002d4",
x"00238",
x"3fc4e",
x"3fce1",
--Row 24
x"00400",
x"00000",
x"3fc00",
x"00000",
x"00400",
x"00000",
x"3fc00",
x"00000",
x"00400",
x"00000",
x"3fc00",
x"00000",
x"00400",
x"00000",
x"3fc00",
x"00000",
x"00400",
x"00000",
x"3fc00",
x"00000",
x"00400",
x"00000",
x"3fc00",
x"00000",
x"00400",
x"00000",
x"3fc00",
x"00000",
x"00400",
x"00000",
x"3fc00",
x"00000",
--Row 25
x"00400",
x"0031f",
x"3fc4e",
x"3fdc8",
x"002d4",
x"00353",
x"3fcf1",
x"3fc14",
x"00000",
x"003ec",
x"0030f",
x"3fcad",
x"3fd2c",
x"00238",
x"003b2",
x"3fce1",
x"3fc00",
x"3fce1",
x"003b2",
x"00238",
x"3fd2c",
x"3fcad",
x"0030f",
x"003ec",
x"00000",
x"3fc14",
x"3fcf1",
x"00353",
x"002d4",
x"3fdc8",
x"3fc4e",
x"0031f",
--Row 26
x"00400",
x"0030f",
x"3fd2c",
x"3fc4e",
x"00000",
x"003b2",
x"002d4",
x"3fcf1",
x"3fc00",
x"3fcf1",
x"002d4",
x"003b2",
x"00000",
x"3fc4e",
x"3fd2c",
x"0030f",
x"00400",
x"0030f",
x"3fd2c",
x"3fc4e",
x"00000",
x"003b2",
x"002d4",
x"3fcf1",
x"3fc00",
x"3fcf1",
x"002d4",
x"003b2",
x"00000",
x"3fc4e",
x"3fd2c",
x"0030f",
--Row 27
x"00400",
x"00238",
x"3fcf1",
x"3fc14",
x"3fd2c",
x"0031f",
x"003b2",
x"00353",
x"00000",
x"3fcad",
x"3fc4e",
x"3fce1",
x"002d4",
x"003ec",
x"0030f",
x"3fdc8",
x"3fc00",
x"3fdc8",
x"0030f",
x"003ec",
x"002d4",
x"3fce1",
x"3fc4e",
x"3fcad",
x"00000",
x"00353",
x"003b2",
x"0031f",
x"3fd2c",
x"3fc14",
x"3fcf1",
x"00238",
--Row 28
x"00400",
x"002d4",
x"00000",
x"3fd2c",
x"3fc00",
x"3fd2c",
x"00000",
x"002d4",
x"00400",
x"002d4",
x"00000",
x"3fd2c",
x"3fc00",
x"3fd2c",
x"00000",
x"002d4",
x"00400",
x"002d4",
x"00000",
x"3fd2c",
x"3fc00",
x"3fd2c",
x"00000",
x"002d4",
x"00400",
x"002d4",
x"00000",
x"3fd2c",
x"3fc00",
x"3fd2c",
x"00000",
x"002d4",
--Row 29
x"00400",
x"00353",
x"0030f",
x"3fce1",
x"3fd2c",
x"3fc14",
x"3fc4e",
x"3fdc8",
x"00000",
x"00238",
x"003b2",
x"003ec",
x"002d4",
x"0031f",
x"3fcf1",
x"3fcad",
x"3fc00",
x"3fcad",
x"3fcf1",
x"0031f",
x"002d4",
x"003ec",
x"003b2",
x"00238",
x"00000",
x"3fdc8",
x"3fc4e",
x"3fc14",
x"3fd2c",
x"3fce1",
x"0030f",
x"00353",
--Row 30
x"00400",
x"003b2",
x"002d4",
x"0030f",
x"00000",
x"3fcf1",
x"3fd2c",
x"3fc4e",
x"3fc00",
x"3fc4e",
x"3fd2c",
x"3fcf1",
x"00000",
x"0030f",
x"002d4",
x"003b2",
x"00400",
x"003b2",
x"002d4",
x"0030f",
x"00000",
x"3fcf1",
x"3fd2c",
x"3fc4e",
x"3fc00",
x"3fc4e",
x"3fd2c",
x"3fcf1",
x"00000",
x"0030f",
x"002d4",
x"003b2",
--Row 31
x"00400",
x"003ec",
x"003b2",
x"00353",
x"002d4",
x"00238",
x"0030f",
x"0031f",
x"00000",
x"3fce1",
x"3fcf1",
x"3fdc8",
x"3fd2c",
x"3fcad",
x"3fc4e",
x"3fc14",
x"3fc00",
x"3fc14",
x"3fc4e",
x"3fcad",
x"3fd2c",
x"3fdc8",
x"3fcf1",
x"3fce1",
x"00000",
x"0031f",
x"0030f",
x"00238",
x"002d4",
x"00353",
x"003b2",
x"003ec"
	
);

BEGIN

	indx <= to_integer(unsigned(index));
	coeff <= memory(indx)(WIDTH-1 downto 0);

END dataflow;
